library verilog;
use verilog.vl_types.all;
entity CODE6C_vlg_vec_tst is
end CODE6C_vlg_vec_tst;
